module manchester_decoder2 (
    input wire aclk,
    input wire aresetn,
    input wire [2:0] bits,
    input wire [2:0] num_bits
);



endmodule
